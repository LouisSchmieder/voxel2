module packet

pub struct ProtocolSettings {
	version int
}
