module read

[id: 0x00]
pub struct StatusRequest {}